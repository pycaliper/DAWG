

`define NUM_WAYS 8
`define NUM_WAYS_WIDTH 3
`define ADDR_WIDTH 32
